//////////////////////////////////////////////////////////////////////////////////
// Company: UW Madison
// Engineer: Jesse Pakula
// 
// Create Date:   
// Design Name: 
// Module Name:    spart 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module spart(
    input clk,
    input rst,
    input iocs,  // I/O chip select, basically enable in this project
    input iorw,	 // I/O Read Not Write bit
    output logic rda,  // receive data available
    output logic tbr,  // transmit buffer ready
    input [1:0] ioaddr,
    inout [7:0] databus,
    output txd,
    input rxd
    );
	
reg [15:0] baud_cnt;
reg [7:0] division_buffer_low;
reg [7:0] division_buffer_high;
reg [15:0] divisor_buffer;
reg [9:0] rx_shift_reg;
reg [9:0] tx_shift_reg;
reg [15:0] rx_middle;
reg [15:0] rx_middle_cnt;
reg [3:0] rx_tx_cnt;
reg [7:0] receive_buffer;
reg [7:0] transmit_buffer;
reg [7:0] status;
reg [7:0] read_data; // multiplexed output of receive buffer and status reg for databus read (ioaddr)
reg [7:0] write_data; // multiplexed output of transmit buffer, DB(Low), and DB(High) based on ioaddr
					 
logic baud_empty;
logic baud_cnt_en;
logic rx_shift_en;
logic tx_shift_en;
logic clr;
logic middle_found; // for checking we are at rxd line
logic rx_middle_en;
logic rx_tx_cnt_en;
logic rx_tx_buf_full;
logic transmit_buffer_en; // enables loading databus into transmission buffer
logic receive_buffer_en;  // enables receiving of data to begin from IO device
logic tx_begin;  // enables loading transmission buffer into tx_shift_reg
logic status_register_read;
logic status_read; // high when reading status register for rda and tbr

logic db_high_en;
logic db_low_en;



// states for SPART
typedef enum reg [3:0] {IDLE, READ, WRITE, RX_FRONT_PORCH, RX, RX_BACK_PORCH, TX_LOAD, TX_FRONT_PORCH, TX, BUFFER_WRITE} state_t;
state_t state, next_state;

// put receive buffer or status reg (depending on ioaddr) on databus if read op
// otherwise high z since SPART will be reading it
assign databus = (iorw) ? read_data : 8'bz;

// first bit of ioaddr is select signal for multiplexer, choosing between status reg and receive_buffer
assign read_data = (ioaddr[0]) ? status : receive_buffer;


// count down divisor buffer
always_ff @(posedge clk, negedge rst) begin
	if (!rst)
		baud_cnt <= divisor_buffer;
	else if (baud_empty)
		baud_cnt <= divisor_buffer;
	else if (baud_cnt_en)
		baud_cnt <= baud_cnt - 16'h0001;  // only count if enable is on
	else
		baud_cnt <= divisor_buffer;	// if we stop counting we want to reset to divisor buffer
end


// status register has rda at bit 0, tbr bit 1, 0s elsewhere.
assign status = {6'b000000, tbr, rda};

// DB_HIGH flop, only load it from data bus when enable signal goes high for 1 clk cycle
always_ff @(posedge clk, negedge rst) begin
	if(!rst)
		// TODO division buffer needs to load starting value based on DIP switches
		division_buffer_high <= 8'b0;
	else if(db_high_en)
		division_buffer_high <= databus;
	else
		division_buffer_high <= division_buffer_high;
end

// DB_LOW flop, only load on enable, otherwise hold value
always_ff @(posedge clk, negedge rst) begin
	if(!rst)
		// TODO load correct starting value based on switches.
		division_buffer_low <= 8'b0;
	else if(db_low_en)
		division_buffer_low <= databus;
	else
		division_buffer_low <= division_buffer_low;
end

// division buffer and baud rate signals
assign baud_empty = (baud_cnt == 16'h0000); // baud_empty when baud_cnt is 0 
assign divisor_buffer = {division_buffer_high[7:0], division_buffer_low[7:0]}; // concatenate for buffer

// TODO find better way to sample in middle of rx line, division is expensive
assign rx_middle = divisor_buffer >> 1'b1; // will sample in middle of bits (divide by 2)

// counter to determine middle_found for correct sampling of rx
always_ff @(posedge clk, negedge rst) begin
	if (!rst)
		rx_middle_cnt <= rx_middle;
	else if (rx_middle_en)
		rx_middle_cnt <= rx_middle_cnt - 16'b1;
	else 
		rx_middle_cnt <= rx_middle; 
end
assign middle_found = (rx_middle_cnt == 0);

// rx and bit counter, include start and stop bits.
always_ff @(posedge clk, negedge rst) begin
	if (!rst)
		rx_tx_cnt <= 4'hA; // always start at 10 for start bit, 8 data, then stop bit
	else if (rx_tx_cnt_en)
		rx_tx_cnt <= rx_tx_cnt - 4'h1; // count down on enable so we know when byte frame ends
	else if (rx_tx_buf_full)
		rx_tx_cnt <= 4'hA; // reload bit counter every time our buffer is full
	else
		rx_tx_cnt <= 4'hA; // reload 10 when enable goes low
end
assign rx_tx_buf_full = (rx_tx_cnt == 4'h0); // signal buffer is full after stop bit
assign rx_tx_cnt_en = rx_shift_en | tx_shift_en; // continue counting when bits are shifted


// rx_shift_reg implementation
always_ff @(posedge clk, negedge rst) begin
	if (!rst)
		rx_shift_reg <= 10'b0;  // 0 on reset
	else if (rx_shift_en)
		rx_shift_reg <= {rxd, rx_shift_reg[9:1]}; // shift rxd from left if enable high
	else 
		rx_shift_reg <= rx_shift_reg; // intentional latch
end

// receive_buffer latches rx_shift data bits when rx_tx_buf_full is asserted
always_ff @(posedge clk, negedge rst) begin
	if (!rst)
		receive_buffer <= 8'b0;
	else if (rx_tx_buf_full)
		receive_buffer <= rx_shift_reg[8:1]; // data bits in middle, start/stop bits on end
	else
		receive_buffer <= receive_buffer; // intentional latch
end

// transmit buffer loads in data from databus when ioaddr enables it
always_ff @(posedge clk, negedge rst) begin
	if (!rst)
		transmit_buffer <= 8'b0;
	else if (transmit_buffer_en)
		transmit_buffer <= databus;  
	else
		transmit_buffer <= transmit_buffer; // intentional latch
end


assign txd = tx_shift_reg[0];  // lsb will be consistently transmitted

// tx_shift_reg implementation
always_ff @(posedge clk, negedge rst) begin
	if (!rst)
		tx_shift_reg <= 10'b1111111111;  // all 1's on reset to hold txd high
	else if(tx_begin)
		tx_shift_reg <= {1'b1, transmit_buffer, 1'b0};
	else if (tx_shift_en)
		tx_shift_reg <= {1'b1, tx_shift_reg[9:1]};
	else
		tx_shift_reg <= tx_shift_reg;  // intentional latch	
end

// rx_shift_en is HIGH in middle of bit being sent: sample in middle of signal
// assign rx_shift_en = middle of bit being sent


// TODO set default signal values
always @(posedge clk, negedge rst) begin
	tbr = 1'b0;
	receive_buffer_en = 1'b0;
	db_high_en = 1'b0;
	db_low_en = 1'b0;
	status_read = 1'b0;
	case(ioaddr)
		2'b00:  
			begin
				if(iorw)
					receive_buffer_en <= 1'b1;
					
				else
					tbr <= 1'b1;
			end
		2'b01:  
			begin
				if(iorw)
					status_read = 1'b1;
				else
					;// nothing
			end
		2'b10:		
			begin
				db_low_en = 1'b1;
			end
		2'b11:
			begin
				db_high_en = 1'b1;
			end
	endcase
end




always_comb begin
	next_state = IDLE; // default state
	rx_middle_en = 1'b0;
	rx_shift_en = 1'b0;
	tx_shift_en = 1'b0;
	tx_begin = 1'b0;
	transmit_buffer_en = 1'b0;
	baud_cnt_en = 1'b0;
	rda = 1'b0;
	
	case(state)
	
		IDLE:
			begin
//				if (iocs & iorw)
//					next_state = READ; NOT SURE IF READ STATE IS NEEDED
				if (iocs & !iorw)
					next_state = WRITE;
				else if (!rxd) // should respond to getting data no matter what, getting data supercedes receiving
					next_state = RX_FRONT_PORCH;
					
				else if (tbr & iocs) // Q: not sure if tbr needs to be a condition here
					next_state = TX_LOAD;
				
				else
					next_state = IDLE;
			end
			
/*		READ:  NOT SURE IF THIS IS NEEDED, THINK IT HAPPENS AUTOMATICALLY
			begin
				
			
			
			end
*/			
		WRITE:
			begin 
				
			
			
			end
			
		RX_FRONT_PORCH:
			begin
				rx_middle_en = 1'b1; // might need to have this in previous state on transition too.
				if (middle_found) begin
					if (!rxd) begin // verify start bit is low
						rx_shift_en = 1'b1;
						next_state = RX; // start sampling data if we have low start bit
					end
					else 
						next_state = IDLE; // back to IDLE if start bit was not low
				end
				else
					next_state = RX_FRONT_PORCH;
			end
		
					
		RX:
			begin
				baud_cnt_en = 1'b1;
				if(baud_empty) begin
					rx_shift_en = 1'b1;
					next_state = RX;
				end
				else if (rx_tx_buf_full) // receive buffer automatically latches on this signal
					if (rx_shift_reg[9]) // check that stop bit was high
						next_state = RX_BACK_PORCH; // done processing this byte
					else
						next_state = IDLE; // go to IDLE if stop bit wasn't high
				else
					next_state = RX;
			end
		
		TX_LOAD:
			begin
				transmit_buffer_en = 1'b1;
				next_state = TX_FRONT_PORCH;
			end
		TX_FRONT_PORCH: 
			begin
				tx_begin = 1'b1;
				next_state = TX;
			end
			
		TX:
			begin
				baud_cnt_en = 1'b1;
				if(baud_empty) begin
					tx_shift_en = 1'b1;
					next_state = TX;
				end
				else if(rx_tx_buf_full)
					next_state = IDLE;
				else
					next_state = TX;
					
			end
			
		// let processor know we have data ready
		RX_BACK_PORCH:
			begin
				rda = 1'b1;
				next_state = IDLE;
			end
			
		
				
	endcase
end

endmodule
